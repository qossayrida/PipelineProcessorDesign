module PipelineProcessor ();
	
	initial begin		 
        #400 $finish; 
    end			
	
	
	
	//******************************************************
	//					clock & registers		
	//******************************************************
	
	wire clk;
	
	
	
	//******************************************************
	//					Control unit registers		
	//****************************************************** 
	
	
	
	
	
	
	//******************************************************
	//					   Pipeline stages		
	//****************************************************** 
	
	
	
endmodule