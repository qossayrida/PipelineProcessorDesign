module PipelineProcessor ();
	

	
	
	
endmodule